RInrery LEGG:
vele IEEE.STO LOGIC 1164.ALL; use IEEE.NOWiRIC TD.ALL:
use IEEE.STOLOGICONSIGNED.ALL;
entity MAIN is
Port (
INPUTS IN STD LOGIc VECTOR r dovnto 0); 
INPVI2 : IN STD:LOGIC—VECTOR r 200.0 0); 
OPR IN STD LOGIC_VECTOR(2 DONNIO 0); 
OVERFLAI OET STD LOGIC;
01 0177 STE_LOGIE_VECTOR (7 elevate 0)
):
end BAIN;
architecture Behavioral of NAIR is
SIGNAL 91 STD_LOGIC:
SIGNAL 92 : STD_LOG/C:
SIGNAL SO : SIM LOGIC;
SIGNAL El : STD_LOGIC_VECTORES DOWNTO 0); SIGNAL 12 STD_LOGIC_VECTOR(2 DOWNTO 0); SIGNAL STD_LOGIC_VECTORI3 WENT ° 0); SIGNAL F2 : STD LOGIC VECTOR13 DGENTO 0); SIGNAL Cl : STDLOGICVECTOR(15 DOMNTO 0); SIGNAL C2 : SIM_LOGIC_VECTOR(IS DM:NW 0); SIGNAL OOTPUT1 SID_LOGIC_VECTOR(15 DONlITO 0); SIGNAL own. STD_LOGIC_VECTOR(31 DOWNTO 0); SIGNAL 091 : STD_LOGIC;
SIGNAL 092 : STD_LOGIC:
SIGNAL 011 SIM_LOGIC_VECTOR(2 DONNED 0); SIGNAL 0E2 : SIT_LOGIC_VECTOR(2 DOWNTO 0); SIGNAL OF1 : STD_LOGIC_VECTOR(9 DUWNTO 0); SIGNAL OF2 : SITLOGICVECTOR(9 DIUNNTO 0);
