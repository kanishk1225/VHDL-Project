LIBRARY IEEE:
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL:
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MAIN is
  Port (
    INPUT1 : IN STD_LOGIC_VECTOR (7 downto 0); 
    INPVI2 : IN STD_LOGIC_VECTOR (7 downto 0); 
    OPR : IN STD_LOGIC_VECTOR (2 downto 0); 
    OVERFLOW : OUT STD_LOGIC;
    01 : OUT STD_LOGIC_VECTOR (7 downto 0)
  ):
end MAIN;

architecture Behavioral of MAIN is

SIGNAL S1 STD_LOGIC:
SIGNAL S2 : STD_LOG/C:
SIGNAL SO : SIM LOGIC;
SIGNAL El : STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL E2 : STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL F1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL F2 : STD LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL Cl : STD_LOGIC_VECTOR(15 DOWNTO 0); 
SIGNAL C2 : STD_LOGIC_VECTOR(IS DOWNTO 0);
SIGNAL OUTPUT1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL OUTPUTX : STD_LOGIC_VECTOR(31 DOWNTO 0); 
SIGNAL OS1 : STD_LOGIC;
SIGNAL OS2 : STD_LOGIC:
SIGNAL OE1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL OE2 : STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL OE1 : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL OF2 : STD_LOGIC_VECTOR(3 DOWNTO 0);

begin
  
MAIN_PROCESS: PROCESS(INPUTI,INPUT2,OPR,E1,FI,C1,E2,F2,C2,OE1,OF1,OE2,OF2,OS1,OS2,OUTPUT1,S1,S2,SO)
BEGIN

OVERFLOW	606:
01 < "0000000n:
51 dcw INPUT1(7);
52 <— INPUT2(7); 
F1(3 DOWNTO 0) <— INPUT1(3 DOWNTO 0);
F2(3 DOWNTO 0) < INPUT 2(3 DOWNTO 0);
E1(2 DOWNTO 0) <— INPUT1(6 DOWNTO 1); 
E2(2 DOWNTO 0) <= INPUT2(6 DOWNTO 4);

IF OUTPUT1(12)='1' THEN
0E1(2 DOWNTO 0)	<- "111";
OF1(3 DOWNTO 0)	<= OUTPUT1(11	TO 8);
ELSIE' OUTPUT1(11)=11' THEN
0E1(2 DOWNTO 0)
